module cpu(
    input             clk,
    input             rst,
    output reg [15:0] addr,
    input      [7:0]  di,
    output reg [7:0]  do,
    output reg        we
);

endmodule
